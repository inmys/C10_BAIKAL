// sopc_top.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module sopc_top (
		input  wire        altpll_0_areset_export,    //   altpll_0_areset.export
		input  wire        altpll_0_inclk0_clk,       //   altpll_0_inclk0.clk
		output wire        altpll_0_locked_export,    //   altpll_0_locked.export
		input  wire        bmc_spi_MISO,              //           bmc_spi.MISO
		output wire        bmc_spi_MOSI,              //                  .MOSI
		output wire        bmc_spi_SCLK,              //                  .SCLK
		output wire        bmc_spi_SS_n,              //                  .SS_n
		input  wire        i2c_0_sda_in,              //             i2c_0.sda_in
		input  wire        i2c_0_scl_in,              //                  .scl_in
		output wire        i2c_0_sda_oe,              //                  .sda_oe
		output wire        i2c_0_scl_oe,              //                  .scl_oe
		input  wire        i2cslave_conduit_data_in,  //          i2cslave.conduit_data_in
		input  wire        i2cslave_conduit_clk_in,   //                  .conduit_clk_in
		output wire        i2cslave_conduit_data_oe,  //                  .conduit_data_oe
		output wire        i2cslave_conduit_clk_oe,   //                  .conduit_clk_oe
		output wire        id32k_clk,                 //             id32k.clk
		input  wire [31:0] pio_in_export,             //            pio_in.export
		output wire [31:0] pio_out_export,            //           pio_out.export
		input  wire        reset_bridge_0_in_reset_n, // reset_bridge_0_in.reset_n
		input  wire        spi_0_MISO,                //             spi_0.MISO
		output wire        spi_0_MOSI,                //                  .MOSI
		output wire        spi_0_SCLK,                //                  .SCLK
		output wire        spi_0_SS_n,                //                  .SS_n
		input  wire        uart_0_sin,                //            uart_0.sin
		output wire        uart_0_sout,               //                  .sout
		output wire        uart_0_sout_oe             //                  .sout_oe
	);

	wire         altpll_0_c0_clk;                                             // altpll_0:c0 -> [a_16550_uart_0:clk, altpll_0:clk, i2c_0:clk, i2cslave_to_avlmm_bridge_0:clk, irq_mapper:clk, jtag_uart_0:clk, mm_bridge_0:clk, mm_interconnect_0:altpll_0_c0_clk, mm_interconnect_1:altpll_0_c0_clk, mm_interconnect_2:altpll_0_c0_clk, nios2_gen2_0:clk, onchip_memory2_0:clk, onchip_memory2_1:clk, onchip_memory2_1:clk2, pio_in:clk, pio_out:clk, rst_controller:clk, spi_0:clk, spi_1:clk, sysid_qsys_0:clock, timer_0:clk]
	wire  [31:0] i2cslave_to_avlmm_bridge_0_avalon_master_readdata;           // mm_interconnect_0:i2cslave_to_avlmm_bridge_0_avalon_master_readdata -> i2cslave_to_avlmm_bridge_0:readdata
	wire         i2cslave_to_avlmm_bridge_0_avalon_master_waitrequest;        // mm_interconnect_0:i2cslave_to_avlmm_bridge_0_avalon_master_waitrequest -> i2cslave_to_avlmm_bridge_0:waitrequest
	wire  [31:0] i2cslave_to_avlmm_bridge_0_avalon_master_address;            // i2cslave_to_avlmm_bridge_0:address -> mm_interconnect_0:i2cslave_to_avlmm_bridge_0_avalon_master_address
	wire         i2cslave_to_avlmm_bridge_0_avalon_master_read;               // i2cslave_to_avlmm_bridge_0:read -> mm_interconnect_0:i2cslave_to_avlmm_bridge_0_avalon_master_read
	wire   [3:0] i2cslave_to_avlmm_bridge_0_avalon_master_byteenable;         // i2cslave_to_avlmm_bridge_0:byteenable -> mm_interconnect_0:i2cslave_to_avlmm_bridge_0_avalon_master_byteenable
	wire         i2cslave_to_avlmm_bridge_0_avalon_master_readdatavalid;      // mm_interconnect_0:i2cslave_to_avlmm_bridge_0_avalon_master_readdatavalid -> i2cslave_to_avlmm_bridge_0:readdatavalid
	wire         i2cslave_to_avlmm_bridge_0_avalon_master_write;              // i2cslave_to_avlmm_bridge_0:write -> mm_interconnect_0:i2cslave_to_avlmm_bridge_0_avalon_master_write
	wire  [31:0] i2cslave_to_avlmm_bridge_0_avalon_master_writedata;          // i2cslave_to_avlmm_bridge_0:writedata -> mm_interconnect_0:i2cslave_to_avlmm_bridge_0_avalon_master_writedata
	wire         mm_interconnect_0_onchip_memory2_1_s1_chipselect;            // mm_interconnect_0:onchip_memory2_1_s1_chipselect -> onchip_memory2_1:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_1_s1_readdata;              // onchip_memory2_1:readdata -> mm_interconnect_0:onchip_memory2_1_s1_readdata
	wire   [5:0] mm_interconnect_0_onchip_memory2_1_s1_address;               // mm_interconnect_0:onchip_memory2_1_s1_address -> onchip_memory2_1:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_1_s1_byteenable;            // mm_interconnect_0:onchip_memory2_1_s1_byteenable -> onchip_memory2_1:byteenable
	wire         mm_interconnect_0_onchip_memory2_1_s1_write;                 // mm_interconnect_0:onchip_memory2_1_s1_write -> onchip_memory2_1:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_1_s1_writedata;             // mm_interconnect_0:onchip_memory2_1_s1_writedata -> onchip_memory2_1:writedata
	wire         mm_interconnect_0_onchip_memory2_1_s1_clken;                 // mm_interconnect_0:onchip_memory2_1_s1_clken -> onchip_memory2_1:clken
	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_1:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_1:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_1:nios2_gen2_0_data_master_debugaccess
	wire  [28:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_1:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_1:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_1:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_1:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_1:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_1:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_1:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [16:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_1:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_1:nios2_gen2_0_instruction_master_read
	wire         nios2_gen2_0_instruction_master_readdatavalid;               // mm_interconnect_1:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire  [31:0] mm_interconnect_1_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_1:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_1_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_1:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_1_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_1_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_1_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_1_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_1_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_1_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_1_altpll_0_pll_slave_readdata;               // altpll_0:readdata -> mm_interconnect_1:altpll_0_pll_slave_readdata
	wire   [1:0] mm_interconnect_1_altpll_0_pll_slave_address;                // mm_interconnect_1:altpll_0_pll_slave_address -> altpll_0:address
	wire         mm_interconnect_1_altpll_0_pll_slave_read;                   // mm_interconnect_1:altpll_0_pll_slave_read -> altpll_0:read
	wire         mm_interconnect_1_altpll_0_pll_slave_write;                  // mm_interconnect_1:altpll_0_pll_slave_write -> altpll_0:write
	wire  [31:0] mm_interconnect_1_altpll_0_pll_slave_writedata;              // mm_interconnect_1:altpll_0_pll_slave_writedata -> altpll_0:writedata
	wire  [31:0] mm_interconnect_1_mm_bridge_0_s0_readdata;                   // mm_bridge_0:s0_readdata -> mm_interconnect_1:mm_bridge_0_s0_readdata
	wire         mm_interconnect_1_mm_bridge_0_s0_waitrequest;                // mm_bridge_0:s0_waitrequest -> mm_interconnect_1:mm_bridge_0_s0_waitrequest
	wire         mm_interconnect_1_mm_bridge_0_s0_debugaccess;                // mm_interconnect_1:mm_bridge_0_s0_debugaccess -> mm_bridge_0:s0_debugaccess
	wire  [11:0] mm_interconnect_1_mm_bridge_0_s0_address;                    // mm_interconnect_1:mm_bridge_0_s0_address -> mm_bridge_0:s0_address
	wire         mm_interconnect_1_mm_bridge_0_s0_read;                       // mm_interconnect_1:mm_bridge_0_s0_read -> mm_bridge_0:s0_read
	wire   [3:0] mm_interconnect_1_mm_bridge_0_s0_byteenable;                 // mm_interconnect_1:mm_bridge_0_s0_byteenable -> mm_bridge_0:s0_byteenable
	wire         mm_interconnect_1_mm_bridge_0_s0_readdatavalid;              // mm_bridge_0:s0_readdatavalid -> mm_interconnect_1:mm_bridge_0_s0_readdatavalid
	wire         mm_interconnect_1_mm_bridge_0_s0_write;                      // mm_interconnect_1:mm_bridge_0_s0_write -> mm_bridge_0:s0_write
	wire  [31:0] mm_interconnect_1_mm_bridge_0_s0_writedata;                  // mm_interconnect_1:mm_bridge_0_s0_writedata -> mm_bridge_0:s0_writedata
	wire   [0:0] mm_interconnect_1_mm_bridge_0_s0_burstcount;                 // mm_interconnect_1:mm_bridge_0_s0_burstcount -> mm_bridge_0:s0_burstcount
	wire         mm_interconnect_1_onchip_memory2_0_s1_chipselect;            // mm_interconnect_1:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_1_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_1:onchip_memory2_0_s1_readdata
	wire  [11:0] mm_interconnect_1_onchip_memory2_0_s1_address;               // mm_interconnect_1:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_1_onchip_memory2_0_s1_byteenable;            // mm_interconnect_1:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_1_onchip_memory2_0_s1_write;                 // mm_interconnect_1:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_1_onchip_memory2_0_s1_writedata;             // mm_interconnect_1:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_1_onchip_memory2_0_s1_clken;                 // mm_interconnect_1:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_bridge_0_m0_waitrequest;                                  // mm_interconnect_2:mm_bridge_0_m0_waitrequest -> mm_bridge_0:m0_waitrequest
	wire  [31:0] mm_bridge_0_m0_readdata;                                     // mm_interconnect_2:mm_bridge_0_m0_readdata -> mm_bridge_0:m0_readdata
	wire         mm_bridge_0_m0_debugaccess;                                  // mm_bridge_0:m0_debugaccess -> mm_interconnect_2:mm_bridge_0_m0_debugaccess
	wire  [11:0] mm_bridge_0_m0_address;                                      // mm_bridge_0:m0_address -> mm_interconnect_2:mm_bridge_0_m0_address
	wire         mm_bridge_0_m0_read;                                         // mm_bridge_0:m0_read -> mm_interconnect_2:mm_bridge_0_m0_read
	wire   [3:0] mm_bridge_0_m0_byteenable;                                   // mm_bridge_0:m0_byteenable -> mm_interconnect_2:mm_bridge_0_m0_byteenable
	wire         mm_bridge_0_m0_readdatavalid;                                // mm_interconnect_2:mm_bridge_0_m0_readdatavalid -> mm_bridge_0:m0_readdatavalid
	wire  [31:0] mm_bridge_0_m0_writedata;                                    // mm_bridge_0:m0_writedata -> mm_interconnect_2:mm_bridge_0_m0_writedata
	wire         mm_bridge_0_m0_write;                                        // mm_bridge_0:m0_write -> mm_interconnect_2:mm_bridge_0_m0_write
	wire   [0:0] mm_bridge_0_m0_burstcount;                                   // mm_bridge_0:m0_burstcount -> mm_interconnect_2:mm_bridge_0_m0_burstcount
	wire         mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_2:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_2:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_2:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_2:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_2:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_2:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_2:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_2_a_16550_uart_0_avalon_slave_readdata;      // a_16550_uart_0:readdata -> mm_interconnect_2:a_16550_uart_0_avalon_slave_readdata
	wire   [8:0] mm_interconnect_2_a_16550_uart_0_avalon_slave_address;       // mm_interconnect_2:a_16550_uart_0_avalon_slave_address -> a_16550_uart_0:addr
	wire         mm_interconnect_2_a_16550_uart_0_avalon_slave_read;          // mm_interconnect_2:a_16550_uart_0_avalon_slave_read -> a_16550_uart_0:read
	wire         mm_interconnect_2_a_16550_uart_0_avalon_slave_write;         // mm_interconnect_2:a_16550_uart_0_avalon_slave_write -> a_16550_uart_0:write
	wire  [31:0] mm_interconnect_2_a_16550_uart_0_avalon_slave_writedata;     // mm_interconnect_2:a_16550_uart_0_avalon_slave_writedata -> a_16550_uart_0:writedata
	wire  [31:0] mm_interconnect_2_sysid_qsys_0_control_slave_readdata;       // sysid_qsys_0:readdata -> mm_interconnect_2:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_2_sysid_qsys_0_control_slave_address;        // mm_interconnect_2:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_2_i2c_0_csr_readdata;                        // i2c_0:readdata -> mm_interconnect_2:i2c_0_csr_readdata
	wire   [3:0] mm_interconnect_2_i2c_0_csr_address;                         // mm_interconnect_2:i2c_0_csr_address -> i2c_0:addr
	wire         mm_interconnect_2_i2c_0_csr_read;                            // mm_interconnect_2:i2c_0_csr_read -> i2c_0:read
	wire         mm_interconnect_2_i2c_0_csr_write;                           // mm_interconnect_2:i2c_0_csr_write -> i2c_0:write
	wire  [31:0] mm_interconnect_2_i2c_0_csr_writedata;                       // mm_interconnect_2:i2c_0_csr_writedata -> i2c_0:writedata
	wire         mm_interconnect_2_pio_out_s1_chipselect;                     // mm_interconnect_2:pio_out_s1_chipselect -> pio_out:chipselect
	wire  [31:0] mm_interconnect_2_pio_out_s1_readdata;                       // pio_out:readdata -> mm_interconnect_2:pio_out_s1_readdata
	wire   [2:0] mm_interconnect_2_pio_out_s1_address;                        // mm_interconnect_2:pio_out_s1_address -> pio_out:address
	wire         mm_interconnect_2_pio_out_s1_write;                          // mm_interconnect_2:pio_out_s1_write -> pio_out:write_n
	wire  [31:0] mm_interconnect_2_pio_out_s1_writedata;                      // mm_interconnect_2:pio_out_s1_writedata -> pio_out:writedata
	wire  [31:0] mm_interconnect_2_pio_in_s1_readdata;                        // pio_in:readdata -> mm_interconnect_2:pio_in_s1_readdata
	wire   [1:0] mm_interconnect_2_pio_in_s1_address;                         // mm_interconnect_2:pio_in_s1_address -> pio_in:address
	wire         mm_interconnect_2_timer_0_s1_chipselect;                     // mm_interconnect_2:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_2_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_2:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_2_timer_0_s1_address;                        // mm_interconnect_2:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_2_timer_0_s1_write;                          // mm_interconnect_2:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_2_timer_0_s1_writedata;                      // mm_interconnect_2:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_2_onchip_memory2_1_s2_chipselect;            // mm_interconnect_2:onchip_memory2_1_s2_chipselect -> onchip_memory2_1:chipselect2
	wire  [31:0] mm_interconnect_2_onchip_memory2_1_s2_readdata;              // onchip_memory2_1:readdata2 -> mm_interconnect_2:onchip_memory2_1_s2_readdata
	wire   [5:0] mm_interconnect_2_onchip_memory2_1_s2_address;               // mm_interconnect_2:onchip_memory2_1_s2_address -> onchip_memory2_1:address2
	wire   [3:0] mm_interconnect_2_onchip_memory2_1_s2_byteenable;            // mm_interconnect_2:onchip_memory2_1_s2_byteenable -> onchip_memory2_1:byteenable2
	wire         mm_interconnect_2_onchip_memory2_1_s2_write;                 // mm_interconnect_2:onchip_memory2_1_s2_write -> onchip_memory2_1:write2
	wire  [31:0] mm_interconnect_2_onchip_memory2_1_s2_writedata;             // mm_interconnect_2:onchip_memory2_1_s2_writedata -> onchip_memory2_1:writedata2
	wire         mm_interconnect_2_onchip_memory2_1_s2_clken;                 // mm_interconnect_2:onchip_memory2_1_s2_clken -> onchip_memory2_1:clken2
	wire         mm_interconnect_2_spi_0_spi_control_port_chipselect;         // mm_interconnect_2:spi_0_spi_control_port_chipselect -> spi_0:spi_select
	wire  [31:0] mm_interconnect_2_spi_0_spi_control_port_readdata;           // spi_0:data_to_cpu -> mm_interconnect_2:spi_0_spi_control_port_readdata
	wire   [2:0] mm_interconnect_2_spi_0_spi_control_port_address;            // mm_interconnect_2:spi_0_spi_control_port_address -> spi_0:mem_addr
	wire         mm_interconnect_2_spi_0_spi_control_port_read;               // mm_interconnect_2:spi_0_spi_control_port_read -> spi_0:read_n
	wire         mm_interconnect_2_spi_0_spi_control_port_write;              // mm_interconnect_2:spi_0_spi_control_port_write -> spi_0:write_n
	wire  [31:0] mm_interconnect_2_spi_0_spi_control_port_writedata;          // mm_interconnect_2:spi_0_spi_control_port_writedata -> spi_0:data_from_cpu
	wire         mm_interconnect_2_spi_1_spi_control_port_chipselect;         // mm_interconnect_2:spi_1_spi_control_port_chipselect -> spi_1:spi_select
	wire  [15:0] mm_interconnect_2_spi_1_spi_control_port_readdata;           // spi_1:data_to_cpu -> mm_interconnect_2:spi_1_spi_control_port_readdata
	wire   [2:0] mm_interconnect_2_spi_1_spi_control_port_address;            // mm_interconnect_2:spi_1_spi_control_port_address -> spi_1:mem_addr
	wire         mm_interconnect_2_spi_1_spi_control_port_read;               // mm_interconnect_2:spi_1_spi_control_port_read -> spi_1:read_n
	wire         mm_interconnect_2_spi_1_spi_control_port_write;              // mm_interconnect_2:spi_1_spi_control_port_write -> spi_1:write_n
	wire  [15:0] mm_interconnect_2_spi_1_spi_control_port_writedata;          // mm_interconnect_2:spi_1_spi_control_port_writedata -> spi_1:data_from_cpu
	wire         irq_mapper_receiver0_irq;                                    // i2c_0:intr -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // timer_0:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                    // spi_0:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                    // spi_1:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                    // a_16550_uart_0:intr -> irq_mapper:receiver5_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [a_16550_uart_0:rst_n, altpll_0:reset, i2c_0:rst_n, i2cslave_to_avlmm_bridge_0:rst_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_bridge_0:reset, mm_interconnect_0:i2cslave_to_avlmm_bridge_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:nios2_gen2_0_reset_reset_bridge_in_reset_reset, mm_interconnect_2:mm_bridge_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory2_0:reset, onchip_memory2_1:reset, onchip_memory2_1:reset2, pio_in:reset_n, pio_out:reset_n, rst_translator:in_reset, spi_0:reset_n, spi_1:reset_n, sysid_qsys_0:reset_n, timer_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, onchip_memory2_1:reset_req, onchip_memory2_1:reset_req2, rst_translator:reset_req_in]

	altera_16550_uart #(
		.FAMILY         ("Cyclone 10 LP"),
		.MEM_BLOCK_TYPE ("AUTO"),
		.FIFO_MODE      (1),
		.FIFO_DEPTH     (256),
		.FIFO_WATERMARK (0),
		.FIFO_HWFC      (1),
		.FIFO_SWFC      (0),
		.DMA_EXTRA      (0)
	) a_16550_uart_0 (
		.addr            (mm_interconnect_2_a_16550_uart_0_avalon_slave_address),   //  avalon_slave.address
		.write           (mm_interconnect_2_a_16550_uart_0_avalon_slave_write),     //              .write
		.writedata       (mm_interconnect_2_a_16550_uart_0_avalon_slave_writedata), //              .writedata
		.read            (mm_interconnect_2_a_16550_uart_0_avalon_slave_read),      //              .read
		.readdata        (mm_interconnect_2_a_16550_uart_0_avalon_slave_readdata),  //              .readdata
		.clk             (altpll_0_c0_clk),                                         //         clock.clk
		.rst_n           (~rst_controller_reset_out_reset),                         //    reset_sink.reset_n
		.intr            (irq_mapper_receiver5_irq),                                //    irq_sender.irq
		.sin             (uart_0_sin),                                              // RS_232_Serial.sin
		.sout            (uart_0_sout),                                             //              .sout
		.sout_oe         (uart_0_sout_oe),                                          //              .sout_oe
		.cts_n           (),                                                        //  RS_232_Modem.cts_n
		.rts_n           (),                                                        //              .rts_n
		.dsr_n           (),                                                        //              .dsr_n
		.dcd_n           (),                                                        //              .dcd_n
		.ri_n            (),                                                        //              .ri_n
		.dtr_n           (),                                                        //              .dtr_n
		.out1_n          (),                                                        //              .out1_n
		.out2_n          (),                                                        //              .out2_n
		.dma_tx_ack_n    (1'b1),                                                    //   (terminated)
		.dma_tx_req_n    (),                                                        //   (terminated)
		.dma_tx_single_n (),                                                        //   (terminated)
		.dma_rx_ack_n    (1'b1),                                                    //   (terminated)
		.dma_rx_req_n    (),                                                        //   (terminated)
		.dma_rx_single_n ()                                                         //   (terminated)
	);

	sopc_top_altpll_0 altpll_0 (
		.clk                (altpll_0_c0_clk),                                //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset),                 // inclk_interface_reset.reset
		.read               (mm_interconnect_1_altpll_0_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_1_altpll_0_pll_slave_write),     //                      .write
		.address            (mm_interconnect_1_altpll_0_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_1_altpll_0_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_1_altpll_0_pll_slave_writedata), //                      .writedata
		.inclk0             (altpll_0_inclk0_clk),                            //                inclk0.clk
		.c0                 (altpll_0_c0_clk),                                //                    c0.clk
		.c1                 (),                                               //                    c1.clk
		.c2                 (id32k_clk),                                      //                    c2.clk
		.areset             (altpll_0_areset_export),                         //        areset_conduit.export
		.locked             (altpll_0_locked_export),                         //        locked_conduit.export
		.scandone           (),                                               //           (terminated)
		.scandataout        (),                                               //           (terminated)
		.phasedone          (),                                               //           (terminated)
		.phasecounterselect (4'b0000),                                        //           (terminated)
		.phaseupdown        (1'b0),                                           //           (terminated)
		.phasestep          (1'b0),                                           //           (terminated)
		.scanclk            (1'b0),                                           //           (terminated)
		.scanclkena         (1'b0),                                           //           (terminated)
		.scandata           (1'b0),                                           //           (terminated)
		.configupdate       (1'b0)                                            //           (terminated)
	);

	altera_avalon_i2c #(
		.USE_AV_ST       (0),
		.FIFO_DEPTH      (64),
		.FIFO_DEPTH_LOG2 (6)
	) i2c_0 (
		.clk       (altpll_0_c0_clk),                       //            clock.clk
		.rst_n     (~rst_controller_reset_out_reset),       //       reset_sink.reset_n
		.intr      (irq_mapper_receiver0_irq),              // interrupt_sender.irq
		.addr      (mm_interconnect_2_i2c_0_csr_address),   //              csr.address
		.read      (mm_interconnect_2_i2c_0_csr_read),      //                 .read
		.write     (mm_interconnect_2_i2c_0_csr_write),     //                 .write
		.writedata (mm_interconnect_2_i2c_0_csr_writedata), //                 .writedata
		.readdata  (mm_interconnect_2_i2c_0_csr_readdata),  //                 .readdata
		.sda_in    (i2c_0_sda_in),                          //       i2c_serial.sda_in
		.scl_in    (i2c_0_scl_in),                          //                 .scl_in
		.sda_oe    (i2c_0_sda_oe),                          //                 .sda_oe
		.scl_oe    (i2c_0_scl_oe),                          //                 .scl_oe
		.src_data  (),                                      //      (terminated)
		.src_valid (),                                      //      (terminated)
		.src_ready (1'b0),                                  //      (terminated)
		.snk_data  (16'b0000000000000000),                  //      (terminated)
		.snk_valid (1'b0),                                  //      (terminated)
		.snk_ready ()                                       //      (terminated)
	);

	altera_i2cslave_to_avlmm_bridge #(
		.I2C_SLAVE_ADDRESS (7'b0100000),
		.BYTE_ADDRESSING   (1),
		.ADDRESS_STEALING  (0),
		.READ_ONLY         (0)
	) i2cslave_to_avlmm_bridge_0 (
		.clk           (altpll_0_c0_clk),                                        //         clock.clk
		.address       (i2cslave_to_avlmm_bridge_0_avalon_master_address),       // avalon_master.address
		.read          (i2cslave_to_avlmm_bridge_0_avalon_master_read),          //              .read
		.readdata      (i2cslave_to_avlmm_bridge_0_avalon_master_readdata),      //              .readdata
		.readdatavalid (i2cslave_to_avlmm_bridge_0_avalon_master_readdatavalid), //              .readdatavalid
		.waitrequest   (i2cslave_to_avlmm_bridge_0_avalon_master_waitrequest),   //              .waitrequest
		.write         (i2cslave_to_avlmm_bridge_0_avalon_master_write),         //              .write
		.byteenable    (i2cslave_to_avlmm_bridge_0_avalon_master_byteenable),    //              .byteenable
		.writedata     (i2cslave_to_avlmm_bridge_0_avalon_master_writedata),     //              .writedata
		.rst_n         (~rst_controller_reset_out_reset),                        //         reset.reset_n
		.i2c_data_in   (i2cslave_conduit_data_in),                               //   conduit_end.conduit_data_in
		.i2c_clk_in    (i2cslave_conduit_clk_in),                                //              .conduit_clk_in
		.i2c_data_oe   (i2cslave_conduit_data_oe),                               //              .conduit_data_oe
		.i2c_clk_oe    (i2cslave_conduit_clk_oe)                                 //              .conduit_clk_oe
	);

	sopc_top_jtag_uart_0 jtag_uart_0 (
		.clk            (altpll_0_c0_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (12),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_0 (
		.clk              (altpll_0_c0_clk),                                //   clk.clk
		.reset            (rst_controller_reset_out_reset),                 // reset.reset
		.s0_waitrequest   (mm_interconnect_1_mm_bridge_0_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_1_mm_bridge_0_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_1_mm_bridge_0_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_1_mm_bridge_0_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_1_mm_bridge_0_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_1_mm_bridge_0_s0_address),       //      .address
		.s0_write         (mm_interconnect_1_mm_bridge_0_s0_write),         //      .write
		.s0_read          (mm_interconnect_1_mm_bridge_0_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_1_mm_bridge_0_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_1_mm_bridge_0_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (mm_bridge_0_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (mm_bridge_0_m0_readdata),                        //      .readdata
		.m0_readdatavalid (mm_bridge_0_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (mm_bridge_0_m0_burstcount),                      //      .burstcount
		.m0_writedata     (mm_bridge_0_m0_writedata),                       //      .writedata
		.m0_address       (mm_bridge_0_m0_address),                         //      .address
		.m0_write         (mm_bridge_0_m0_write),                           //      .write
		.m0_read          (mm_bridge_0_m0_read),                            //      .read
		.m0_byteenable    (mm_bridge_0_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (mm_bridge_0_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                               // (terminated)
		.m0_response      (2'b00)                                           // (terminated)
	);

	sopc_top_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (altpll_0_c0_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                           //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	sopc_top_onchip_memory2_0 onchip_memory2_0 (
		.clk        (altpll_0_c0_clk),                                  //   clk1.clk
		.address    (mm_interconnect_1_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_1_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_1_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_1_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_1_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_1_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_1_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	sopc_top_onchip_memory2_1 onchip_memory2_1 (
		.clk         (altpll_0_c0_clk),                                  //   clk1.clk
		.address     (mm_interconnect_0_onchip_memory2_1_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_onchip_memory2_1_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_onchip_memory2_1_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_onchip_memory2_1_s1_write),      //       .write
		.readdata    (mm_interconnect_0_onchip_memory2_1_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_onchip_memory2_1_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_onchip_memory2_1_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),               //       .reset_req
		.address2    (mm_interconnect_2_onchip_memory2_1_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_2_onchip_memory2_1_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_2_onchip_memory2_1_s2_clken),      //       .clken
		.write2      (mm_interconnect_2_onchip_memory2_1_s2_write),      //       .write
		.readdata2   (mm_interconnect_2_onchip_memory2_1_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_2_onchip_memory2_1_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_2_onchip_memory2_1_s2_byteenable), //       .byteenable
		.clk2        (altpll_0_c0_clk),                                  //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),                   // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze      (1'b0)                                              // (terminated)
	);

	sopc_top_pio_in pio_in (
		.clk      (altpll_0_c0_clk),                      //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_2_pio_in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_2_pio_in_s1_readdata), //                    .readdata
		.in_port  (pio_in_export)                         // external_connection.export
	);

	sopc_top_pio_out pio_out (
		.clk        (altpll_0_c0_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_2_pio_out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_pio_out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_pio_out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_pio_out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_pio_out_s1_readdata),   //                    .readdata
		.out_port   (pio_out_export)                           // external_connection.export
	);

	sopc_top_spi_0 spi_0 (
		.clk           (altpll_0_c0_clk),                                     //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                     //            reset.reset_n
		.data_from_cpu (mm_interconnect_2_spi_0_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_2_spi_0_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_2_spi_0_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_2_spi_0_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_2_spi_0_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_2_spi_0_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver3_irq),                            //              irq.irq
		.MISO          (spi_0_MISO),                                          //         external.export
		.MOSI          (spi_0_MOSI),                                          //                 .export
		.SCLK          (spi_0_SCLK),                                          //                 .export
		.SS_n          (spi_0_SS_n)                                           //                 .export
	);

	sopc_top_spi_1 spi_1 (
		.clk           (altpll_0_c0_clk),                                     //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                     //            reset.reset_n
		.data_from_cpu (mm_interconnect_2_spi_1_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_2_spi_1_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_2_spi_1_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_2_spi_1_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_2_spi_1_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_2_spi_1_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver4_irq),                            //              irq.irq
		.MISO          (bmc_spi_MISO),                                        //         external.export
		.MOSI          (bmc_spi_MOSI),                                        //                 .export
		.SCLK          (bmc_spi_SCLK),                                        //                 .export
		.SS_n          (bmc_spi_SS_n)                                         //                 .export
	);

	sopc_top_sysid_qsys_0 sysid_qsys_0 (
		.clock    (altpll_0_c0_clk),                                       //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_2_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_2_sysid_qsys_0_control_slave_address)   //              .address
	);

	sopc_top_timer_0 timer_0 (
		.clk        (altpll_0_c0_clk),                         //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_2_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_2_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_2_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_2_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_2_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                 //   irq.irq
	);

	sopc_top_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c0_clk                                              (altpll_0_c0_clk),                                        //                                            altpll_0_c0.clk
		.i2cslave_to_avlmm_bridge_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                         // i2cslave_to_avlmm_bridge_0_reset_reset_bridge_in_reset.reset
		.i2cslave_to_avlmm_bridge_0_avalon_master_address             (i2cslave_to_avlmm_bridge_0_avalon_master_address),       //               i2cslave_to_avlmm_bridge_0_avalon_master.address
		.i2cslave_to_avlmm_bridge_0_avalon_master_waitrequest         (i2cslave_to_avlmm_bridge_0_avalon_master_waitrequest),   //                                                       .waitrequest
		.i2cslave_to_avlmm_bridge_0_avalon_master_byteenable          (i2cslave_to_avlmm_bridge_0_avalon_master_byteenable),    //                                                       .byteenable
		.i2cslave_to_avlmm_bridge_0_avalon_master_read                (i2cslave_to_avlmm_bridge_0_avalon_master_read),          //                                                       .read
		.i2cslave_to_avlmm_bridge_0_avalon_master_readdata            (i2cslave_to_avlmm_bridge_0_avalon_master_readdata),      //                                                       .readdata
		.i2cslave_to_avlmm_bridge_0_avalon_master_readdatavalid       (i2cslave_to_avlmm_bridge_0_avalon_master_readdatavalid), //                                                       .readdatavalid
		.i2cslave_to_avlmm_bridge_0_avalon_master_write               (i2cslave_to_avlmm_bridge_0_avalon_master_write),         //                                                       .write
		.i2cslave_to_avlmm_bridge_0_avalon_master_writedata           (i2cslave_to_avlmm_bridge_0_avalon_master_writedata),     //                                                       .writedata
		.onchip_memory2_1_s1_address                                  (mm_interconnect_0_onchip_memory2_1_s1_address),          //                                    onchip_memory2_1_s1.address
		.onchip_memory2_1_s1_write                                    (mm_interconnect_0_onchip_memory2_1_s1_write),            //                                                       .write
		.onchip_memory2_1_s1_readdata                                 (mm_interconnect_0_onchip_memory2_1_s1_readdata),         //                                                       .readdata
		.onchip_memory2_1_s1_writedata                                (mm_interconnect_0_onchip_memory2_1_s1_writedata),        //                                                       .writedata
		.onchip_memory2_1_s1_byteenable                               (mm_interconnect_0_onchip_memory2_1_s1_byteenable),       //                                                       .byteenable
		.onchip_memory2_1_s1_chipselect                               (mm_interconnect_0_onchip_memory2_1_s1_chipselect),       //                                                       .chipselect
		.onchip_memory2_1_s1_clken                                    (mm_interconnect_0_onchip_memory2_1_s1_clken)             //                                                       .clken
	);

	sopc_top_mm_interconnect_1 mm_interconnect_1 (
		.altpll_0_c0_clk                                (altpll_0_c0_clk),                                            //                              altpll_0_c0.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                             // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                           //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                       //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                        //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                              //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                          //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                             //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                         //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                       //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                    //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                       //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                   //                                         .readdata
		.nios2_gen2_0_instruction_master_readdatavalid  (nios2_gen2_0_instruction_master_readdatavalid),              //                                         .readdatavalid
		.altpll_0_pll_slave_address                     (mm_interconnect_1_altpll_0_pll_slave_address),               //                       altpll_0_pll_slave.address
		.altpll_0_pll_slave_write                       (mm_interconnect_1_altpll_0_pll_slave_write),                 //                                         .write
		.altpll_0_pll_slave_read                        (mm_interconnect_1_altpll_0_pll_slave_read),                  //                                         .read
		.altpll_0_pll_slave_readdata                    (mm_interconnect_1_altpll_0_pll_slave_readdata),              //                                         .readdata
		.altpll_0_pll_slave_writedata                   (mm_interconnect_1_altpll_0_pll_slave_writedata),             //                                         .writedata
		.mm_bridge_0_s0_address                         (mm_interconnect_1_mm_bridge_0_s0_address),                   //                           mm_bridge_0_s0.address
		.mm_bridge_0_s0_write                           (mm_interconnect_1_mm_bridge_0_s0_write),                     //                                         .write
		.mm_bridge_0_s0_read                            (mm_interconnect_1_mm_bridge_0_s0_read),                      //                                         .read
		.mm_bridge_0_s0_readdata                        (mm_interconnect_1_mm_bridge_0_s0_readdata),                  //                                         .readdata
		.mm_bridge_0_s0_writedata                       (mm_interconnect_1_mm_bridge_0_s0_writedata),                 //                                         .writedata
		.mm_bridge_0_s0_burstcount                      (mm_interconnect_1_mm_bridge_0_s0_burstcount),                //                                         .burstcount
		.mm_bridge_0_s0_byteenable                      (mm_interconnect_1_mm_bridge_0_s0_byteenable),                //                                         .byteenable
		.mm_bridge_0_s0_readdatavalid                   (mm_interconnect_1_mm_bridge_0_s0_readdatavalid),             //                                         .readdatavalid
		.mm_bridge_0_s0_waitrequest                     (mm_interconnect_1_mm_bridge_0_s0_waitrequest),               //                                         .waitrequest
		.mm_bridge_0_s0_debugaccess                     (mm_interconnect_1_mm_bridge_0_s0_debugaccess),               //                                         .debugaccess
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_address),     //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_write),       //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_read),        //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_readdata),    //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_writedata),   //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_byteenable),  //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_waitrequest), //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_debugaccess), //                                         .debugaccess
		.onchip_memory2_0_s1_address                    (mm_interconnect_1_onchip_memory2_0_s1_address),              //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_1_onchip_memory2_0_s1_write),                //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_1_onchip_memory2_0_s1_readdata),             //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_1_onchip_memory2_0_s1_writedata),            //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_1_onchip_memory2_0_s1_byteenable),           //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_1_onchip_memory2_0_s1_chipselect),           //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_1_onchip_memory2_0_s1_clken)                 //                                         .clken
	);

	sopc_top_mm_interconnect_2 mm_interconnect_2 (
		.altpll_0_c0_clk                               (altpll_0_c0_clk),                                             //                             altpll_0_c0.clk
		.mm_bridge_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // mm_bridge_0_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_m0_address                        (mm_bridge_0_m0_address),                                      //                          mm_bridge_0_m0.address
		.mm_bridge_0_m0_waitrequest                    (mm_bridge_0_m0_waitrequest),                                  //                                        .waitrequest
		.mm_bridge_0_m0_burstcount                     (mm_bridge_0_m0_burstcount),                                   //                                        .burstcount
		.mm_bridge_0_m0_byteenable                     (mm_bridge_0_m0_byteenable),                                   //                                        .byteenable
		.mm_bridge_0_m0_read                           (mm_bridge_0_m0_read),                                         //                                        .read
		.mm_bridge_0_m0_readdata                       (mm_bridge_0_m0_readdata),                                     //                                        .readdata
		.mm_bridge_0_m0_readdatavalid                  (mm_bridge_0_m0_readdatavalid),                                //                                        .readdatavalid
		.mm_bridge_0_m0_write                          (mm_bridge_0_m0_write),                                        //                                        .write
		.mm_bridge_0_m0_writedata                      (mm_bridge_0_m0_writedata),                                    //                                        .writedata
		.mm_bridge_0_m0_debugaccess                    (mm_bridge_0_m0_debugaccess),                                  //                                        .debugaccess
		.a_16550_uart_0_avalon_slave_address           (mm_interconnect_2_a_16550_uart_0_avalon_slave_address),       //             a_16550_uart_0_avalon_slave.address
		.a_16550_uart_0_avalon_slave_write             (mm_interconnect_2_a_16550_uart_0_avalon_slave_write),         //                                        .write
		.a_16550_uart_0_avalon_slave_read              (mm_interconnect_2_a_16550_uart_0_avalon_slave_read),          //                                        .read
		.a_16550_uart_0_avalon_slave_readdata          (mm_interconnect_2_a_16550_uart_0_avalon_slave_readdata),      //                                        .readdata
		.a_16550_uart_0_avalon_slave_writedata         (mm_interconnect_2_a_16550_uart_0_avalon_slave_writedata),     //                                        .writedata
		.i2c_0_csr_address                             (mm_interconnect_2_i2c_0_csr_address),                         //                               i2c_0_csr.address
		.i2c_0_csr_write                               (mm_interconnect_2_i2c_0_csr_write),                           //                                        .write
		.i2c_0_csr_read                                (mm_interconnect_2_i2c_0_csr_read),                            //                                        .read
		.i2c_0_csr_readdata                            (mm_interconnect_2_i2c_0_csr_readdata),                        //                                        .readdata
		.i2c_0_csr_writedata                           (mm_interconnect_2_i2c_0_csr_writedata),                       //                                        .writedata
		.jtag_uart_0_avalon_jtag_slave_address         (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_address),     //           jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write           (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_write),       //                                        .write
		.jtag_uart_0_avalon_jtag_slave_read            (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_read),        //                                        .read
		.jtag_uart_0_avalon_jtag_slave_readdata        (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_readdata),    //                                        .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata       (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_writedata),   //                                        .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest     (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                        .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect      (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                        .chipselect
		.onchip_memory2_1_s2_address                   (mm_interconnect_2_onchip_memory2_1_s2_address),               //                     onchip_memory2_1_s2.address
		.onchip_memory2_1_s2_write                     (mm_interconnect_2_onchip_memory2_1_s2_write),                 //                                        .write
		.onchip_memory2_1_s2_readdata                  (mm_interconnect_2_onchip_memory2_1_s2_readdata),              //                                        .readdata
		.onchip_memory2_1_s2_writedata                 (mm_interconnect_2_onchip_memory2_1_s2_writedata),             //                                        .writedata
		.onchip_memory2_1_s2_byteenable                (mm_interconnect_2_onchip_memory2_1_s2_byteenable),            //                                        .byteenable
		.onchip_memory2_1_s2_chipselect                (mm_interconnect_2_onchip_memory2_1_s2_chipselect),            //                                        .chipselect
		.onchip_memory2_1_s2_clken                     (mm_interconnect_2_onchip_memory2_1_s2_clken),                 //                                        .clken
		.pio_in_s1_address                             (mm_interconnect_2_pio_in_s1_address),                         //                               pio_in_s1.address
		.pio_in_s1_readdata                            (mm_interconnect_2_pio_in_s1_readdata),                        //                                        .readdata
		.pio_out_s1_address                            (mm_interconnect_2_pio_out_s1_address),                        //                              pio_out_s1.address
		.pio_out_s1_write                              (mm_interconnect_2_pio_out_s1_write),                          //                                        .write
		.pio_out_s1_readdata                           (mm_interconnect_2_pio_out_s1_readdata),                       //                                        .readdata
		.pio_out_s1_writedata                          (mm_interconnect_2_pio_out_s1_writedata),                      //                                        .writedata
		.pio_out_s1_chipselect                         (mm_interconnect_2_pio_out_s1_chipselect),                     //                                        .chipselect
		.spi_0_spi_control_port_address                (mm_interconnect_2_spi_0_spi_control_port_address),            //                  spi_0_spi_control_port.address
		.spi_0_spi_control_port_write                  (mm_interconnect_2_spi_0_spi_control_port_write),              //                                        .write
		.spi_0_spi_control_port_read                   (mm_interconnect_2_spi_0_spi_control_port_read),               //                                        .read
		.spi_0_spi_control_port_readdata               (mm_interconnect_2_spi_0_spi_control_port_readdata),           //                                        .readdata
		.spi_0_spi_control_port_writedata              (mm_interconnect_2_spi_0_spi_control_port_writedata),          //                                        .writedata
		.spi_0_spi_control_port_chipselect             (mm_interconnect_2_spi_0_spi_control_port_chipselect),         //                                        .chipselect
		.spi_1_spi_control_port_address                (mm_interconnect_2_spi_1_spi_control_port_address),            //                  spi_1_spi_control_port.address
		.spi_1_spi_control_port_write                  (mm_interconnect_2_spi_1_spi_control_port_write),              //                                        .write
		.spi_1_spi_control_port_read                   (mm_interconnect_2_spi_1_spi_control_port_read),               //                                        .read
		.spi_1_spi_control_port_readdata               (mm_interconnect_2_spi_1_spi_control_port_readdata),           //                                        .readdata
		.spi_1_spi_control_port_writedata              (mm_interconnect_2_spi_1_spi_control_port_writedata),          //                                        .writedata
		.spi_1_spi_control_port_chipselect             (mm_interconnect_2_spi_1_spi_control_port_chipselect),         //                                        .chipselect
		.sysid_qsys_0_control_slave_address            (mm_interconnect_2_sysid_qsys_0_control_slave_address),        //              sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata           (mm_interconnect_2_sysid_qsys_0_control_slave_readdata),       //                                        .readdata
		.timer_0_s1_address                            (mm_interconnect_2_timer_0_s1_address),                        //                              timer_0_s1.address
		.timer_0_s1_write                              (mm_interconnect_2_timer_0_s1_write),                          //                                        .write
		.timer_0_s1_readdata                           (mm_interconnect_2_timer_0_s1_readdata),                       //                                        .readdata
		.timer_0_s1_writedata                          (mm_interconnect_2_timer_0_s1_writedata),                      //                                        .writedata
		.timer_0_s1_chipselect                         (mm_interconnect_2_timer_0_s1_chipselect)                      //                                        .chipselect
	);

	sopc_top_irq_mapper irq_mapper (
		.clk           (altpll_0_c0_clk),                //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_bridge_0_in_reset_n),         // reset_in0.reset
		.clk            (altpll_0_c0_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
